module uart_reg_tb;
    reg clk = 0; rst = 0;
    reg wr_i, rd_i;
    reg rx_fifo_empty_i;
    reg [7:0] rx_fifo_in;
    reg [2:0] addr_i;
    reg [7:0] din_i;
    reg rx_oe, rx_pe, rx_fe, rx_bi;
    wire tx_push_o; //add new data to Tx fifo
    wire rx_pop_o; //read data from Rx fifo

    wire baud_out;

    wire tx_rst, rx_rst;
    wire [3:0] rx_fifo_threshold;
 
    wire [7:0] dout_o;
 
    csr_t csr;

    regs_uart dut (
                    .clk(clk),
                    .rst(rst),
                    .wr_i(wr_i),
                    .rd_i(rd_i),
                    .rx_fifo_empty_i(rx_fifo_empty_i),
                    .rx_oe(rx_oe),
                    .rx_pe(rx_pe),
                    .rx_fe(rx_fe),
                    .rx_bi(rx_bi),
                    .addr_i(addr_i),
                    .din_i(din_i),
                    .tx_push_o(tx_push_o),
                    .rx_pop_o(rx_pop_o),
                    .baud_out(baud_out),
                    .tx_rst(tx_rst),
                    .rx_rst(rx_rst),
                    .rx_fifo_threshold(rx_fifo_threshold),
                    .dout_o(dout_o),
                    .csr(csr),
                    .rx_fifo_in(rx_fifo_in)
                    
    );

    always #5 clk = ~clk;

    initial begin
        rst = 1;
        repeat(5) @(posedge clk);
        rst = 0;
        /////// update lsb and msb of divisor
        //////// sel DLAB(msb) of lcr (3H) reg to 1
        @(negedge clk);
        wr_i = 1;
        addr_i = 3'h3;
        din_i <= 8'1000_0000;

       /////////////// Update LSB of divisor latch
       @(negedge clk);
       addr_i = 3'h0;
       din_i <= 8'b0000_1000; //08


       //////////// Update MSB of divisor latch
       @(negedge clk)
       addr_i = 3'h1;
       din_i <= 8'b0000_00001;

       //////////////Make DLAB 0 
       @(negedge clk)
       addr_i = 3'h3;
       din_i <= 8'b0000_00000;
       $finish; 
    end

    
endmodule